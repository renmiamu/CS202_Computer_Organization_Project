module ALU (
    input [3:0] ALUop,
    input [31:0] ALU_input_1,
    input [31:0] ALU_input_2,
    
);
    
endmodule