module IO (
    
);
    
endmodule