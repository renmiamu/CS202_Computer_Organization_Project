module swtich (
    input clk,
    input rst
    
);
    
endmodule